library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity instruction_memory is										
port ( i_ADDR : in  std_logic_vector(31 downto 0);  -- Endereço de memória
       o_OUT  : out std_logic_vector(31 downto 0)); -- Dados de saída
end instruction_memory;
	
architecture arq_1 of instruction_memory is
  type t_MEMORY is array (0 to 255) of std_logic_vector (31 downto 0); -- Cria um tipo memory_array que e um vetor de 256 posicoes que guarda 32 bits em cada uma delas
  signal w_MEM : t_MEMORY := (
    0  => "00000000000000000000010000010011",
    1  => "00000000000000000000010010010011",
    2  => "00000000000100000000101010010011",
    3  => "00000000010100000000100100010011",
    4  => "00000000100101001000001010110011",
    5  => "00000000010100101000001010110011",
    6  => "00000000010101000000001010110011",
    7  => "00000001001000101010000000100011",
    8  => "00000001010101001010001010110011",
    9  => "00000010000000101000111001100011",
    10 => "00000001010101001000010010110011",
    11 => "01000001010110010000100100110011",
    12 => "00000000100101001000001010110011",
    13 => "00000000010100101000001010110011",
    14 => "00000000010101000000001010110011",
    15 => "00000001001000101010000000100011",
    16 => "00000001010101001010001010110011",
    17 => "00000000000000101000111001100011",
    18 => "00000001010101001000010010110011",
    19 => "01000001010110010000100100110011",
    20 => "00000000100101001000001010110011",
    21 => "00000000010100101000001010110011",
    22 => "00000000010101000000001010110011",
    23 => "00000001001000101010000000100011",
    24 => "00000000100101001000001010110011",
    25 => "00000000010100101000001010110011",
    26 => "00000000010101000000001010110011",
    27 => "00000000000000101010001100000011",
    28 => "01000001010101001000010010110011",
    29 => "00000000100101001000001010110011",
    30 => "00000000010100101000001010110011",
    31 => "00000000010101000000001010110011",
    32 => "00000000000000101010001110000011",
    33 => "00000000011100110000111000110011",
    34 => "00000000000000000000000000010011",
    others => (others => '0')
  );
	
begin 
  o_OUT <= w_MEM(to_integer(unsigned(i_ADDR(9 downto 2))));
end arq_1;